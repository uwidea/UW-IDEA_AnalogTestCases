** Generated for: hspiceD
** Generated on: Jan  5 07:55:36 2020
** Design library name: AP_SerDes
** Design cell name: Bias_v2
** Design view name: schematic
.PARAM w3 w4 w1mn w w2p w1m w3p


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65LP/models/hspice/toplevel.l" tt_lib

** Library name: AP_SerDes
** Cell name: Bias_v2
** View name: schematic
m24<19> in_1m net0159 net0136<0> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<18> in_1m net0159 net0136<1> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<17> in_1m net0159 net0136<2> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<16> in_1m net0159 net0136<3> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<15> in_1m net0159 net0136<4> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<14> in_1m net0159 net0136<5> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<13> in_1m net0159 net0136<6> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<12> in_1m net0159 net0136<7> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<11> in_1m net0159 net0136<8> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<10> in_1m net0159 net0136<9> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m29<9> net0184<0> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<8> net0184<1> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<7> net0184<2> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<6> net0184<3> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m27<0> net073 net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m26<5> net0220<0> net0159 net0165<0> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<4> net0220<1> net0159 net0165<1> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<3> net0220<2> net0159 net0165<2> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m25<9> net0162<0> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<8> net0162<1> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<7> net0162<2> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<6> net0162<3> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m23<0> net081 net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m29<5> net0187<0> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<4> net0187<1> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<3> net0187<2> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m28<0> net0228 net0159 net073 avss nch l=1e-6 w='w3*1' m=100 nf=1 
m24<2> net0232<0> net0159 net0154<0> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<1> net0232<1> net0159 net0154<1> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m28<2> net0200<0> net0159 net0179<0> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<1> net0200<1> net0159 net0179<1> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m95<5> in_5m calin5<2> net0196<0> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m95<4> in_5m calin5<2> net0196<1> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m95<3> in_5m calin5<2> net0196<2> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m24<5> net0227<0> net0159 net0145<0> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<4> net0227<1> net0159 net0145<1> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<3> net0227<2> net0159 net0145<2> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m23<9> net0140<0> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<8> net0140<1> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<7> net0140<2> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<6> net0140<3> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m27<9> net0173<0> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<8> net0173<1> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<7> net0173<2> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<6> net0173<3> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m25<0> net077 net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m100<5> in_7m calin7<2> net0210<0> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m100<4> in_7m calin7<2> net0210<1> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m100<3> in_7m calin7<2> net0210<2> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m99<2> in_7m calin7<1> net0214<0> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m99<1> in_7m calin7<1> net0214<1> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m98<0> in_7m calin7<0> net062 avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m97<0> in_5m calin5<0> net0228 avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m30<0> net062 net0159 net069 avss nch l=1e-6 w='w3*1' m=140 nf=1 
m23<5> net0145<0> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<4> net0145<1> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<3> net0145<2> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m96<2> in_5m calin5<1> net0200<0> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m96<1> in_5m calin5<1> net0200<1> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m93<9> in_3m calin3<3> net0178<0> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m93<8> in_3m calin3<3> net0178<1> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m93<7> in_3m calin3<3> net0178<2> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m93<6> in_3m calin3<3> net0178<3> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m94<9> in_5m calin5<3> net0192<0> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m94<8> in_5m calin5<3> net0192<1> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m94<7> in_5m calin5<3> net0192<2> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m94<6> in_5m calin5<3> net0192<3> avss nch l=250e-9 w='w1mn*1' m=100 nf=1 
m25<5> net0165<0> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<4> net0165<1> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<3> net0165<2> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m74<9> in_1m calin1<3> net0157<0> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m74<8> in_1m calin1<3> net0157<1> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m74<7> in_1m calin1<3> net0157<2> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m74<6> in_1m calin1<3> net0157<3> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m90<0> in_3m calin3<0> net078 avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m30<19> in_7m net0159 net0182<0> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<18> in_7m net0159 net0182<1> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<17> in_7m net0159 net0182<2> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<16> in_7m net0159 net0182<3> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<15> in_7m net0159 net0182<4> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<14> in_7m net0159 net0182<5> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<13> in_7m net0159 net0182<6> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<12> in_7m net0159 net0182<7> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<11> in_7m net0159 net0182<8> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<10> in_7m net0159 net0182<9> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m91<2> in_3m calin3<1> net0186<0> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m91<1> in_3m calin3<1> net0186<1> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m30<5> net0210<0> net0159 net0187<0> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<4> net0210<1> net0159 net0187<1> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<3> net0210<2> net0159 net0187<2> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m28<19> in_5m net0159 net0171<0> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<18> in_5m net0159 net0171<1> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<17> in_5m net0159 net0171<2> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<16> in_5m net0159 net0171<3> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<15> in_5m net0159 net0171<4> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<14> in_5m net0159 net0171<5> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<13> in_5m net0159 net0171<6> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<12> in_5m net0159 net0171<7> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<11> in_5m net0159 net0171<8> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<10> in_5m net0159 net0171<9> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<5> net0196<0> net0159 net0176<0> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<4> net0196<1> net0159 net0176<1> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<3> net0196<2> net0159 net0176<2> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m26<19> in_3m net0159 net0160<0> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<18> in_3m net0159 net0160<1> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<17> in_3m net0159 net0160<2> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<16> in_3m net0159 net0160<3> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<15> in_3m net0159 net0160<4> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<14> in_3m net0159 net0160<5> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<13> in_3m net0159 net0160<6> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<12> in_3m net0159 net0160<7> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<11> in_3m net0159 net0160<8> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<10> in_3m net0159 net0160<9> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m92<5> in_3m calin3<2> net0220<0> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m92<4> in_3m calin3<2> net0220<1> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m92<3> in_3m calin3<2> net0220<2> avss nch l=250e-9 w='w1mn*1' m=60 nf=1 
m29<0> net069 net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m23<2> net0154<0> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<1> net0154<1> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m30<2> net0214<0> net0159 net0190<0> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<1> net0214<1> net0159 net0190<1> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m27<2> net0179<0> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<1> net0179<1> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m101<9> in_7m calin7<3> net0206<0> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m101<8> in_7m calin7<3> net0206<1> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m101<7> in_7m calin7<3> net0206<2> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m101<6> in_7m calin7<3> net0206<3> avss nch l=250e-9 w='w1mn*1' m=140 nf=1 
m26<2> net0186<0> net0159 net0168<0> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<1> net0186<1> net0159 net0168<1> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m27<5> net0176<0> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<4> net0176<1> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<3> net0176<2> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m26<0> net078 net0159 net077 avss nch l=1e-6 w='w3*1' m=60 nf=1 
m24<0> net0222 net0159 net081 avss nch l=1e-6 w='w3*1' m=20 nf=1 
m102<5> in_1m calin1<2> net0227<0> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m102<4> in_1m calin1<2> net0227<1> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m102<3> in_1m calin1<2> net0227<2> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m25<2> net0168<0> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<1> net0168<1> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m104<0> in_1m calin1<0> net0222 avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m29<2> net0190<0> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<1> net0190<1> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m103<2> in_1m calin1<1> net0232<0> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m103<1> in_1m calin1<1> net0232<1> avss nch l=250e-9 w='w1mn*1' m=20 nf=1 
m30<9> net0206<0> net0159 net0184<0> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<8> net0206<1> net0159 net0184<1> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<7> net0206<2> net0159 net0184<2> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m30<6> net0206<3> net0159 net0184<3> avss nch l=1e-6 w='w3*1' m=140 nf=1 
m28<9> net0192<0> net0159 net0173<0> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<8> net0192<1> net0159 net0173<1> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<7> net0192<2> net0159 net0173<2> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m28<6> net0192<3> net0159 net0173<3> avss nch l=1e-6 w='w3*1' m=100 nf=1 
m29<19> net0182<0> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<18> net0182<1> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<17> net0182<2> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<16> net0182<3> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<15> net0182<4> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<14> net0182<5> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<13> net0182<6> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<12> net0182<7> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<11> net0182<8> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m29<10> net0182<9> net0159 avss avss nch l=1e-6 w='w4*1' m=140 nf=1 
m26<9> net0178<0> net0159 net0162<0> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<8> net0178<1> net0159 net0162<1> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<7> net0178<2> net0159 net0162<2> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m26<6> net0178<3> net0159 net0162<3> avss nch l=1e-6 w='w3*1' m=60 nf=1 
m27<19> net0171<0> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<18> net0171<1> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<17> net0171<2> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<16> net0171<3> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<15> net0171<4> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<14> net0171<5> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<13> net0171<6> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<12> net0171<7> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<11> net0171<8> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m27<10> net0171<9> net0159 avss avss nch l=1e-6 w='w4*1' m=100 nf=1 
m24<9> net0157<0> net0159 net0140<0> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<8> net0157<1> net0159 net0140<1> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<7> net0157<2> net0159 net0140<2> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m24<6> net0157<3> net0159 net0140<3> avss nch l=1e-6 w='w3*1' m=20 nf=1 
m25<19> net0160<0> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<18> net0160<1> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<17> net0160<2> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<16> net0160<3> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<15> net0160<4> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<14> net0160<5> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<13> net0160<6> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<12> net0160<7> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<11> net0160<8> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m25<10> net0160<9> net0159 avss avss nch l=1e-6 w='w4*1' m=60 nf=1 
m13<19> net0159 net0159 net067<0> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<18> net0159 net0159 net067<1> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<17> net0159 net0159 net067<2> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<16> net0159 net0159 net067<3> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<15> net0159 net0159 net067<4> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<14> net0159 net0159 net067<5> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<13> net0159 net0159 net067<6> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<12> net0159 net0159 net067<7> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<11> net0159 net0159 net067<8> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<10> net0159 net0159 net067<9> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<9> net0159 net0159 net067<10> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<8> net0159 net0159 net067<11> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<7> net0159 net0159 net067<12> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<6> net0159 net0159 net067<13> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<5> net0159 net0159 net067<14> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<4> net0159 net0159 net067<15> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<3> net0159 net0159 net067<16> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<2> net0159 net0159 net067<17> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<1> net0159 net0159 net067<18> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m13<0> net0159 net0159 net067<19> avss nch l=1e-6 w='w3*1' m=1 nf=1 
m23<19> net0136<0> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<18> net0136<1> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<17> net0136<2> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<16> net0136<3> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<15> net0136<4> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<14> net0136<5> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<13> net0136<6> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<12> net0136<7> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<11> net0136<8> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m23<10> net0136<9> net0159 avss avss nch l=1e-6 w='w4*1' m=20 nf=1 
m14<19> net067<0> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<18> net067<1> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<17> net067<2> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<16> net067<3> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<15> net067<4> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<14> net067<5> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<13> net067<6> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<12> net067<7> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<11> net067<8> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<10> net067<9> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<9> net067<10> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<8> net067<11> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<7> net067<12> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<6> net067<13> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<5> net067<14> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<4> net067<15> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<3> net067<16> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<2> net067<17> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<1> net067<18> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m14<0> net067<19> net0159 avss avss nch l=1e-6 w='w4*1' m=1 nf=1 
m4 net011 ibg avss avss nch l=2e-6 w='w*1' m=1 nf=1 
m3 ibg ibg avss avss nch l=2e-6 w='w*1' m=1 nf=1 
m33<9> net0163<0> net011 net089<0> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<8> net0163<1> net011 net089<1> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<7> net0163<2> net011 net089<2> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<6> net0163<3> net011 net089<3> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m82<2> ip_5m calip5<1> net0180<0> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m82<1> ip_5m calip5<1> net0180<1> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m31<0> net0107 net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m33<2> net0169<0> net011 net091<0> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<1> net0169<1> net011 net091<1> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m86<5> ip_7m calip7<2> net0188<0> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m86<4> ip_7m calip7<2> net0188<1> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m86<3> ip_7m calip7<2> net0188<2> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m85<2> ip_7m calip7<1> net0191<0> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m85<1> ip_7m calip7<1> net0191<1> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m84<0> ip_7m calip7<0> net057 avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m83<0> ip_5m calip5<0> net0195 avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m38<0> net041 net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m31<5> net085<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<4> net085<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<3> net085<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m37<2> net0191<0> net011 net0101<0> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<1> net0191<1> net011 net0101<1> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m36<5> net0177<0> net011 net096<0> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<4> net0177<1> net011 net096<1> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<3> net0177<2> net011 net096<2> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m87<9> ip_7m calip7<3> net0185<0> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m87<8> ip_7m calip7<3> net0185<1> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m87<7> ip_7m calip7<3> net0185<2> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m87<6> ip_7m calip7<3> net0185<3> avdd pch l=100e-9 w='w1m*1' m=140 nf=1 
m32<2> net0113<0> net011 net086<0> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<1> net0113<1> net011 net086<1> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m81<5> ip_5m calip5<2> net0177<0> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m81<4> ip_5m calip5<2> net0177<1> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m81<3> ip_5m calip5<2> net0177<2> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m80<9> ip_5m calip5<3> net0174<0> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m80<8> ip_5m calip5<3> net0174<1> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m80<7> ip_5m calip5<3> net0174<2> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m80<6> ip_5m calip5<3> net0174<3> avdd pch l=100e-9 w='w1m*1' m=100 nf=1 
m79<9> ip_3m calip3<3> net0163<0> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m79<8> ip_3m calip3<3> net0163<1> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m79<7> ip_3m calip3<3> net0163<2> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m79<6> ip_3m calip3<3> net0163<3> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m36<9> net0174<0> net011 net095<0> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<8> net0174<1> net011 net095<1> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<7> net0174<2> net011 net095<2> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<6> net0174<3> net011 net095<3> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m78<5> ip_3m calip3<2> net0166<0> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m78<4> ip_3m calip3<2> net0166<1> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m78<3> ip_3m calip3<2> net0166<2> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m37<0> net057 net011 net041 avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m32<0> net0117 net011 net0107 avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m35<5> net096<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<4> net096<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<3> net096<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m33<0> net033 net011 net0105 avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m31<2> net086<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<1> net086<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m36<2> net0180<0> net011 net097<0> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<1> net0180<1> net011 net097<1> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m34<2> net091<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<1> net091<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m31<9> net084<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<8> net084<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<7> net084<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<6> net084<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m35<2> net097<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<1> net097<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m34<0> net0105 net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m38<2> net0101<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<1> net0101<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m32<5> net0125<0> net011 net085<0> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<4> net0125<1> net011 net085<1> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<3> net0125<2> net011 net085<2> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m37<5> net0188<0> net011 net0100<0> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<4> net0188<1> net011 net0100<1> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<3> net0188<2> net011 net0100<2> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m35<0> net0106 net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m33<5> net0166<0> net011 net090<0> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<4> net0166<1> net011 net090<1> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<3> net0166<2> net011 net090<2> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m32<9> net0124<0> net011 net084<0> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<8> net0124<1> net011 net084<1> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<7> net0124<2> net011 net084<2> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<6> net0124<3> net011 net084<3> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m35<19> net093<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<18> net093<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<17> net093<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<16> net093<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<15> net093<4> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<14> net093<5> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<13> net093<6> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<12> net093<7> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<11> net093<8> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<10> net093<9> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m31<19> net083<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<18> net083<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<17> net083<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<16> net083<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<15> net083<4> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<14> net083<5> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<13> net083<6> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<12> net083<7> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<11> net083<8> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m31<10> net083<9> net011 avdd avdd pch l=1e-6 w='w3p*1' m=20 nf=1 
m72<9> ip_1m calip1<3> net0124<0> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<8> ip_1m calip1<3> net0124<1> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<7> ip_1m calip1<3> net0124<2> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<6> ip_1m calip1<3> net0124<3> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m76<0> ip_3m calip3<0> net033 avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m72<0> ip_1m calip1<0> net0117 avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<2> ip_1m calip1<1> net0113<0> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<1> ip_1m calip1<1> net0113<1> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<5> ip_1m calip1<2> net0125<0> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<4> ip_1m calip1<2> net0125<1> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m72<3> ip_1m calip1<2> net0125<2> avdd pch l=100e-9 w='w1m*1' m=20 nf=1 
m38<19> net098<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<18> net098<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<17> net098<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<16> net098<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<15> net098<4> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<14> net098<5> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<13> net098<6> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<12> net098<7> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<11> net098<8> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<10> net098<9> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m77<2> ip_3m calip3<1> net0169<0> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m77<1> ip_3m calip3<1> net0169<1> avdd pch l=100e-9 w='w1m*1' m=60 nf=1 
m37<9> net0185<0> net011 net099<0> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<8> net0185<1> net011 net099<1> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<7> net0185<2> net011 net099<2> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<6> net0185<3> net011 net099<3> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m36<0> net0195 net011 net0106 avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m38<5> net0100<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<4> net0100<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<3> net0100<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m34<19> net088<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<18> net088<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<17> net088<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<16> net088<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<15> net088<4> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<14> net088<5> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<13> net088<6> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<12> net088<7> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<11> net088<8> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<10> net088<9> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m38<9> net099<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<8> net099<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<7> net099<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m38<6> net099<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=140 nf=1 
m37<19> ip_7m net011 net098<0> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<18> ip_7m net011 net098<1> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<17> ip_7m net011 net098<2> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<16> ip_7m net011 net098<3> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<15> ip_7m net011 net098<4> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<14> ip_7m net011 net098<5> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<13> ip_7m net011 net098<6> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<12> ip_7m net011 net098<7> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<11> ip_7m net011 net098<8> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m37<10> ip_7m net011 net098<9> avdd pch l=1e-6 w='w2p*1' m=140 nf=1 
m35<9> net095<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<8> net095<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<7> net095<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m35<6> net095<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=100 nf=1 
m34<9> net089<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<8> net089<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<7> net089<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<6> net089<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m36<19> ip_5m net011 net093<0> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<18> ip_5m net011 net093<1> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<17> ip_5m net011 net093<2> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<16> ip_5m net011 net093<3> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<15> ip_5m net011 net093<4> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<14> ip_5m net011 net093<5> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<13> ip_5m net011 net093<6> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<12> ip_5m net011 net093<7> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<11> ip_5m net011 net093<8> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m36<10> ip_5m net011 net093<9> avdd pch l=1e-6 w='w2p*1' m=100 nf=1 
m33<19> ip_3m net011 net088<0> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<18> ip_3m net011 net088<1> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<17> ip_3m net011 net088<2> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<16> ip_3m net011 net088<3> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<15> ip_3m net011 net088<4> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<14> ip_3m net011 net088<5> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<13> ip_3m net011 net088<6> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<12> ip_3m net011 net088<7> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<11> ip_3m net011 net088<8> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m33<10> ip_3m net011 net088<9> avdd pch l=1e-6 w='w2p*1' m=60 nf=1 
m34<5> net090<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<4> net090<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m34<3> net090<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=60 nf=1 
m32<19> ip_1m net011 net083<0> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<18> ip_1m net011 net083<1> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<17> ip_1m net011 net083<2> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<16> ip_1m net011 net083<3> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<15> ip_1m net011 net083<4> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<14> ip_1m net011 net083<5> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<13> ip_1m net011 net083<6> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<12> ip_1m net011 net083<7> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<11> ip_1m net011 net083<8> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m32<10> ip_1m net011 net083<9> avdd pch l=1e-6 w='w2p*1' m=20 nf=1 
m10<19> net0159 net011 net046<0> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<18> net0159 net011 net046<1> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<17> net0159 net011 net046<2> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<16> net0159 net011 net046<3> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<15> net0159 net011 net046<4> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<14> net0159 net011 net046<5> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<13> net0159 net011 net046<6> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<12> net0159 net011 net046<7> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<11> net0159 net011 net046<8> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<10> net0159 net011 net046<9> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<9> net0159 net011 net046<10> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<8> net0159 net011 net046<11> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<7> net0159 net011 net046<12> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<6> net0159 net011 net046<13> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<5> net0159 net011 net046<14> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<4> net0159 net011 net046<15> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<3> net0159 net011 net046<16> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<2> net0159 net011 net046<17> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<1> net0159 net011 net046<18> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m10<0> net0159 net011 net046<19> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<19> net011 net011 net045<0> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<18> net011 net011 net045<1> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<17> net011 net011 net045<2> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<16> net011 net011 net045<3> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<15> net011 net011 net045<4> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<14> net011 net011 net045<5> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<13> net011 net011 net045<6> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<12> net011 net011 net045<7> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<11> net011 net011 net045<8> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<10> net011 net011 net045<9> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<9> net011 net011 net045<10> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<8> net011 net011 net045<11> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<7> net011 net011 net045<12> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<6> net011 net011 net045<13> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<5> net011 net011 net045<14> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<4> net011 net011 net045<15> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<3> net011 net011 net045<16> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<2> net011 net011 net045<17> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<1> net011 net011 net045<18> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m7<0> net011 net011 net045<19> avdd pch l=1e-6 w='w2p*1' m=1 nf=1 
m9<19> net046<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<18> net046<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<17> net046<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<16> net046<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<15> net046<4> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<14> net046<5> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<13> net046<6> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<12> net046<7> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<11> net046<8> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<10> net046<9> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<9> net046<10> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<8> net046<11> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<7> net046<12> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<6> net046<13> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<5> net046<14> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<4> net046<15> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<3> net046<16> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<2> net046<17> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<1> net046<18> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m9<0> net046<19> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<19> net045<0> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<18> net045<1> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<17> net045<2> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<16> net045<3> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<15> net045<4> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<14> net045<5> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<13> net045<6> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<12> net045<7> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<11> net045<8> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<10> net045<9> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<9> net045<10> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<8> net045<11> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<7> net045<12> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<6> net045<13> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<5> net045<14> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<4> net045<15> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<3> net045<16> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<2> net045<17> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<1> net045<18> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
m8<0> net045<19> net011 avdd avdd pch l=1e-6 w='w3p*1' m=1 nf=1 
.END

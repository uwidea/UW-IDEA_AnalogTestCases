** Generated for: hspiceD
** Generated on: Jan  5 03:09:29 2020
** Design library name: civicR
** Design cell name: DLDO_TOP
** Design view name: schematic


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/home/lab.apps/vlsiapps/kits/tsmc/N65LP/models/hspice/toplevel.l" tt_lib

** Library name: tcbn65lp
** Cell name: DFQD1
** View name: schematic
.subckt DFQD1 d cp q vdd vss
m0 net7 net13 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi4 net24 net63 vss vss nch l=60e-9 w=370e-9 m=1 nf=1 
mi56 net37 net7 vss vss nch l=60e-9 w=150e-9 m=1 nf=1 
m1 net11 net67 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi50 net11 net25 net13 vss nch l=60e-9 w=190e-9 m=1 nf=1 
m2 net25 net63 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi5 net67 d net24 vss nch l=60e-9 w=370e-9 m=1 nf=1 
m3 net63 cp vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi49 net13 net63 net37 vss nch l=60e-9 w=150e-9 m=1 nf=1 
mi48 net9 net11 vss vss nch l=60e-9 w=150e-9 m=1 nf=1 
m4 q net7 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi47 net67 net25 net9 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m5 net7 net13 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m6 net25 net63 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi43 net56 net11 vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi6 net67 d net49 vdd pch l=60e-9 w=460e-9 m=1 nf=1 
m7 net63 cp vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m8 q net7 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi57 net13 net25 net72 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
m9 net11 net67 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi52 net11 net63 net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi51 net72 net7 vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi45 net67 net63 net56 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi7 net49 net25 vdd vdd pch l=60e-9 w=460e-9 m=1 nf=1 
.ends DFQD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: INVD1
** View name: schematic
.subckt INVD1 i zn vdd vss
m0 zn i vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 zn i vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends INVD1
** End of subcircuit definition.

** Library name: civic
** Cell name: ULDO4HVT
** View name: schematic
.subckt ULDO4HVT a d en rs vdd vo vss z
m16 vss vo vss vss nch_hvt l=130e-9 w=795e-9 m=1 nf=1 
m18 z rs net027 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m0 net027 net020 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m14 net021 en vss vss nch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m13 net21 d net021 vss nch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m20 net020 a vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m10 vo net21 vdd vdd pch_hvt l=60e-9 w=1.88e-6 m=1 nf=1 
m1 z rs vo vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m15 net21 en vdd vdd pch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m12 net21 d vdd vdd pch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m19 net020 a vo vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m17 z net020 vo vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends ULDO4HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: DCAP16HVT
** View name: schematic
.subckt DCAP16HVT vdd vss
mi4 vss net11 vss vss nch_hvt l=690e-9 w=300e-9 m=1 nf=1 
mi8 vss net11 vss vss nch_hvt l=690e-9 w=300e-9 m=1 nf=1 
m_u2 net5 net11 vss vss nch_hvt l=60e-9 w=300e-9 m=1 nf=1 
mi7 vss net11 vss vss nch_hvt l=690e-9 w=300e-9 m=1 nf=1 
mi3 vdd net5 vdd vdd pch_hvt l=690e-9 w=430e-9 m=1 nf=1 
mi6 vdd net5 vdd vdd pch_hvt l=690e-9 w=430e-9 m=1 nf=1 
m_u1 net11 net5 vdd vdd pch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi5 vdd net5 vdd vdd pch_hvt l=690e-9 w=430e-9 m=1 nf=1 
.ends DCAP16HVT
** End of subcircuit definition.

** Library name: civic
** Cell name: ULDO_BANK
** View name: schematic
.subckt ULDO_BANK code<5> code<4> code<3> code<2> code<1> code<0> en ro<0> ro<64> ro<63> ro<62> ro<61> ro<60> ro<59> ro<58> ro<57> ro<56> ro<55> ro<54> ro<53> ro<52> ro<51> ro<50> ro<49> ro<48> ro<47> ro<46> ro<45> ro<44> ro<43> ro<42> ro<41> ro<40> ro<39> ro<38> ro<37> ro<36> ro<35> ro<34> ro<33> ro<32> ro<31> ro<30> ro<29> ro<28> ro<27> ro<26> ro<25> ro<24> ro<23> ro<22> ro<21> ro<20> ro<19> ro<18> ro<17> ro<16> ro<15> ro<14> ro<13> ro<12> ro<11> ro<10> ro<9> ro<8> ro<7> ro<6> ro<5> ro<4> ro<3> ro<2> ro<1> rs_rising vdd vout vss
xpwb14<3> ro<44> code<4> en rs_rising vdd vout vss ro<45> ULDO4HVT
xpwb14<2> ro<45> code<4> en rs_rising vdd vout vss ro<46> ULDO4HVT
xpwb14<1> ro<46> code<3> en rs_rising vdd vout vss ro<47> ULDO4HVT
xpwb14<0> ro<47> code<3> en rs_rising vdd vout vss ro<48> ULDO4HVT
xpwb7<3> ro<28> code<4> en rs_rising vdd vout vss ro<29> ULDO4HVT
xpwb7<2> ro<29> code<4> en rs_rising vdd vout vss ro<30> ULDO4HVT
xpwb7<1> ro<30> code<2> en rs_rising vdd vout vss ro<31> ULDO4HVT
xpwb7<0> ro<31> code<2> en rs_rising vdd vout vss ro<32> ULDO4HVT
xpwb6<3> ro<12> code<5> en rs_rising vdd vout vss ro<13> ULDO4HVT
xpwb6<2> ro<13> code<5> en rs_rising vdd vout vss ro<14> ULDO4HVT
xpwb6<1> ro<14> code<5> en rs_rising vdd vout vss ro<15> ULDO4HVT
xpwb6<0> ro<15> code<5> en rs_rising vdd vout vss ro<16> ULDO4HVT
xpwb15<3> ro<60> code<4> en rs_rising vdd vout vss ro<61> ULDO4HVT
xpwb15<2> ro<61> code<4> en rs_rising vdd vout vss ro<62> ULDO4HVT
xpwb15<1> ro<62> code<3> en rs_rising vdd vout vss ro<63> ULDO4HVT
xpwb15<0> ro<63> code<3> en rs_rising vdd vout vss ro<64> ULDO4HVT
xpwb13<3> ro<56> code<4> en rs_rising vdd vout vss ro<57> ULDO4HVT
xpwb13<2> ro<57> code<4> en rs_rising vdd vout vss ro<58> ULDO4HVT
xpwb13<1> ro<58> code<3> en rs_rising vdd vout vss ro<59> ULDO4HVT
xpwb13<0> ro<59> code<3> en rs_rising vdd vout vss ro<60> ULDO4HVT
xpwb12<3> ro<40> code<5> en rs_rising vdd vout vss ro<41> ULDO4HVT
xpwb12<2> ro<41> code<5> en rs_rising vdd vout vss ro<42> ULDO4HVT
xpwb12<1> ro<42> code<5> en rs_rising vdd vout vss ro<43> ULDO4HVT
xpwb12<0> ro<43> code<1> en rs_rising vdd vout vss ro<44> ULDO4HVT
xpwb5<3> ro<24> code<5> en rs_rising vdd vout vss ro<25> ULDO4HVT
xpwb5<2> ro<25> code<5> en rs_rising vdd vout vss ro<26> ULDO4HVT
xpwb5<1> ro<26> code<5> en rs_rising vdd vout vss ro<27> ULDO4HVT
xpwb5<0> ro<27> code<0> en rs_rising vdd vout vss ro<28> ULDO4HVT
xpwb4<3> ro<8> code<5> en rs_rising vdd vout vss ro<9> ULDO4HVT
xpwb4<2> ro<9> code<5> en rs_rising vdd vout vss ro<10> ULDO4HVT
xpwb4<1> ro<10> code<5> en rs_rising vdd vout vss ro<11> ULDO4HVT
xpwb4<0> ro<11> code<5> en rs_rising vdd vout vss ro<12> ULDO4HVT
xpwb11<3> ro<52> code<5> en rs_rising vdd vout vss ro<53> ULDO4HVT
xpwb11<2> ro<53> code<5> en rs_rising vdd vout vss ro<54> ULDO4HVT
xpwb11<1> ro<54> code<3> en rs_rising vdd vout vss ro<55> ULDO4HVT
xpwb11<0> ro<55> code<3> en rs_rising vdd vout vss ro<56> ULDO4HVT
xpwb10<3> ro<36> code<5> en rs_rising vdd vout vss ro<37> ULDO4HVT
xpwb10<2> ro<37> code<5> en rs_rising vdd vout vss ro<38> ULDO4HVT
xpwb10<1> ro<38> code<5> en rs_rising vdd vout vss ro<39> ULDO4HVT
xpwb10<0> ro<39> code<1> en rs_rising vdd vout vss ro<40> ULDO4HVT
xpwb3<3> ro<20> code<5> en rs_rising vdd vout vss ro<21> ULDO4HVT
xpwb3<2> ro<21> code<5> en rs_rising vdd vout vss ro<22> ULDO4HVT
xpwb3<1> ro<22> code<2> en rs_rising vdd vout vss ro<23> ULDO4HVT
xpwb3<0> ro<23> code<2> en rs_rising vdd vout vss ro<24> ULDO4HVT
xpwb2<3> ro<4> code<5> en rs_rising vdd vout vss ro<5> ULDO4HVT
xpwb2<2> ro<5> code<5> en rs_rising vdd vout vss ro<6> ULDO4HVT
xpwb2<1> ro<6> code<5> en rs_rising vdd vout vss ro<7> ULDO4HVT
xpwb2<0> ro<7> code<5> en rs_rising vdd vout vss ro<8> ULDO4HVT
xpwb9<3> ro<48> code<4> en rs_rising vdd vout vss ro<49> ULDO4HVT
xpwb9<2> ro<49> code<4> en rs_rising vdd vout vss ro<50> ULDO4HVT
xpwb9<1> ro<50> code<4> en rs_rising vdd vout vss ro<51> ULDO4HVT
xpwb9<0> ro<51> code<4> en rs_rising vdd vout vss ro<52> ULDO4HVT
xpbw8<3> ro<32> code<5> en rs_rising vdd vout vss ro<33> ULDO4HVT
xpbw8<2> ro<33> code<5> en rs_rising vdd vout vss ro<34> ULDO4HVT
xpbw8<1> ro<34> code<5> en rs_rising vdd vout vss ro<35> ULDO4HVT
xpbw8<0> ro<35> code<5> en rs_rising vdd vout vss ro<36> ULDO4HVT
xpwb1<3> ro<16> code<4> en rs_rising vdd vout vss ro<17> ULDO4HVT
xpwb1<2> ro<17> code<4> en rs_rising vdd vout vss ro<18> ULDO4HVT
xpwb1<1> ro<18> code<4> en rs_rising vdd vout vss ro<19> ULDO4HVT
xpwb1<0> ro<19> code<4> en rs_rising vdd vout vss ro<20> ULDO4HVT
xpwb0<3> ro<0> code<5> en rs_rising vdd vout vss ro<1> ULDO4HVT
xpwb0<2> ro<1> code<5> en rs_rising vdd vout vss ro<2> ULDO4HVT
xpwb0<1> ro<2> code<5> en rs_rising vdd vout vss ro<3> ULDO4HVT
xpwb0<0> ro<3> en en rs_rising vdd vout vss ro<4> ULDO4HVT
xddcp<47> vdd vss DCAP16HVT
xddcp<46> vdd vss DCAP16HVT
xddcp<45> vdd vss DCAP16HVT
xddcp<44> vdd vss DCAP16HVT
xddcp<43> vdd vss DCAP16HVT
xddcp<42> vdd vss DCAP16HVT
xddcp<41> vdd vss DCAP16HVT
xddcp<40> vdd vss DCAP16HVT
xddcp<39> vdd vss DCAP16HVT
xddcp<38> vdd vss DCAP16HVT
xddcp<37> vdd vss DCAP16HVT
xddcp<36> vdd vss DCAP16HVT
xddcp<35> vdd vss DCAP16HVT
xddcp<34> vdd vss DCAP16HVT
xddcp<33> vdd vss DCAP16HVT
xddcp<32> vdd vss DCAP16HVT
xddcp<31> vdd vss DCAP16HVT
xddcp<30> vdd vss DCAP16HVT
xddcp<29> vdd vss DCAP16HVT
xddcp<28> vdd vss DCAP16HVT
xddcp<27> vdd vss DCAP16HVT
xddcp<26> vdd vss DCAP16HVT
xddcp<25> vdd vss DCAP16HVT
xddcp<24> vdd vss DCAP16HVT
xddcp<23> vdd vss DCAP16HVT
xddcp<22> vdd vss DCAP16HVT
xddcp<21> vdd vss DCAP16HVT
xddcp<20> vdd vss DCAP16HVT
xddcp<19> vdd vss DCAP16HVT
xddcp<18> vdd vss DCAP16HVT
xddcp<17> vdd vss DCAP16HVT
xddcp<16> vdd vss DCAP16HVT
xddcp<15> vdd vss DCAP16HVT
xddcp<14> vdd vss DCAP16HVT
xddcp<13> vdd vss DCAP16HVT
xddcp<12> vdd vss DCAP16HVT
xddcp<11> vdd vss DCAP16HVT
xddcp<10> vdd vss DCAP16HVT
xddcp<9> vdd vss DCAP16HVT
xddcp<8> vdd vss DCAP16HVT
xddcp<7> vdd vss DCAP16HVT
xddcp<6> vdd vss DCAP16HVT
xddcp<5> vdd vss DCAP16HVT
xddcp<4> vdd vss DCAP16HVT
xddcp<3> vdd vss DCAP16HVT
xddcp<2> vdd vss DCAP16HVT
xddcp<1> vdd vss DCAP16HVT
xddcp<0> vdd vss DCAP16HVT
.ends ULDO_BANK
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: INVD0HVT
** View name: schematic
.subckt INVD0HVT i zn vdd vss
m0 zn i vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m1 zn i vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
.ends INVD0HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: ND2D0HVT
** View name: schematic
.subckt ND2D0HVT a1 a2 zn vdd vss
m0 zn a1 net1 vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m1 net1 a2 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m2 zn a1 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
m3 zn a2 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
.ends ND2D0HVT
** End of subcircuit definition.

** Library name: civic
** Cell name: Dlvlxft_16B
** View name: schematic
.subckt Dlvlxft_16B bus_in<15> bus_in<14> bus_in<13> bus_in<12> bus_in<11> bus_in<10> bus_in<9> bus_in<8> bus_in<7> bus_in<6> bus_in<5> bus_in<4> bus_in<3> bus_in<2> bus_in<1> bus_in<0> bus_out<15> bus_out<14> bus_out<13> bus_out<12> bus_out<11> bus_out<10> bus_out<9> bus_out<8> bus_out<7> bus_out<6> bus_out<5> bus_out<4> bus_out<3> bus_out<2> bus_out<1> bus_out<0> bus_outn<15> bus_outn<14> bus_outn<13> bus_outn<12> bus_outn<11> bus_outn<10> bus_outn<9> bus_outn<8> bus_outn<7> bus_outn<6> bus_outn<5> bus_outn<4> bus_outn<3> bus_outn<2> bus_outn<1> bus_outn<0> vdd vss
xi2<15> bus_in<15> n<15> vdd vss INVD0HVT
xi2<14> bus_in<14> n<14> vdd vss INVD0HVT
xi2<13> bus_in<13> n<13> vdd vss INVD0HVT
xi2<12> bus_in<12> n<12> vdd vss INVD0HVT
xi2<11> bus_in<11> n<11> vdd vss INVD0HVT
xi2<10> bus_in<10> n<10> vdd vss INVD0HVT
xi2<9> bus_in<9> n<9> vdd vss INVD0HVT
xi2<8> bus_in<8> n<8> vdd vss INVD0HVT
xi2<7> bus_in<7> n<7> vdd vss INVD0HVT
xi2<6> bus_in<6> n<6> vdd vss INVD0HVT
xi2<5> bus_in<5> n<5> vdd vss INVD0HVT
xi2<4> bus_in<4> n<4> vdd vss INVD0HVT
xi2<3> bus_in<3> n<3> vdd vss INVD0HVT
xi2<2> bus_in<2> n<2> vdd vss INVD0HVT
xi2<1> bus_in<1> n<1> vdd vss INVD0HVT
xi2<0> bus_in<0> n<0> vdd vss INVD0HVT
xi1<15> n<15> bus_outn<15> bus_out<15> vdd vss ND2D0HVT
xi1<14> n<14> bus_outn<14> bus_out<14> vdd vss ND2D0HVT
xi1<13> n<13> bus_outn<13> bus_out<13> vdd vss ND2D0HVT
xi1<12> n<12> bus_outn<12> bus_out<12> vdd vss ND2D0HVT
xi1<11> n<11> bus_outn<11> bus_out<11> vdd vss ND2D0HVT
xi1<10> n<10> bus_outn<10> bus_out<10> vdd vss ND2D0HVT
xi1<9> n<9> bus_outn<9> bus_out<9> vdd vss ND2D0HVT
xi1<8> n<8> bus_outn<8> bus_out<8> vdd vss ND2D0HVT
xi1<7> n<7> bus_outn<7> bus_out<7> vdd vss ND2D0HVT
xi1<6> n<6> bus_outn<6> bus_out<6> vdd vss ND2D0HVT
xi1<5> n<5> bus_outn<5> bus_out<5> vdd vss ND2D0HVT
xi1<4> n<4> bus_outn<4> bus_out<4> vdd vss ND2D0HVT
xi1<3> n<3> bus_outn<3> bus_out<3> vdd vss ND2D0HVT
xi1<2> n<2> bus_outn<2> bus_out<2> vdd vss ND2D0HVT
xi1<1> n<1> bus_outn<1> bus_out<1> vdd vss ND2D0HVT
xi1<0> n<0> bus_outn<0> bus_out<0> vdd vss ND2D0HVT
xi3<15> bus_in<15> bus_out<15> bus_outn<15> vdd vss ND2D0HVT
xi3<14> bus_in<14> bus_out<14> bus_outn<14> vdd vss ND2D0HVT
xi3<13> bus_in<13> bus_out<13> bus_outn<13> vdd vss ND2D0HVT
xi3<12> bus_in<12> bus_out<12> bus_outn<12> vdd vss ND2D0HVT
xi3<11> bus_in<11> bus_out<11> bus_outn<11> vdd vss ND2D0HVT
xi3<10> bus_in<10> bus_out<10> bus_outn<10> vdd vss ND2D0HVT
xi3<9> bus_in<9> bus_out<9> bus_outn<9> vdd vss ND2D0HVT
xi3<8> bus_in<8> bus_out<8> bus_outn<8> vdd vss ND2D0HVT
xi3<7> bus_in<7> bus_out<7> bus_outn<7> vdd vss ND2D0HVT
xi3<6> bus_in<6> bus_out<6> bus_outn<6> vdd vss ND2D0HVT
xi3<5> bus_in<5> bus_out<5> bus_outn<5> vdd vss ND2D0HVT
xi3<4> bus_in<4> bus_out<4> bus_outn<4> vdd vss ND2D0HVT
xi3<3> bus_in<3> bus_out<3> bus_outn<3> vdd vss ND2D0HVT
xi3<2> bus_in<2> bus_out<2> bus_outn<2> vdd vss ND2D0HVT
xi3<1> bus_in<1> bus_out<1> bus_outn<1> vdd vss ND2D0HVT
xi3<0> bus_in<0> bus_out<0> bus_outn<0> vdd vss ND2D0HVT
.ends Dlvlxft_16B
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: CKND1HVT
** View name: schematic
.subckt CKND1HVT i zn vdd vss
m_u2 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u1 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends CKND1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: MUX3D1HVT
** View name: schematic
.subckt MUX3D1HVT i0 i1 i2 s0 s1 z vdd vss
m0 net37 net13 net25 vss nch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m1 net33 s0 net25 vss nch_hvt l=60e-9 w=240e-9 m=1 nf=1 
m2 net37 i0 vss vss nch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m3 net25 net9 net79 vss nch_hvt l=60e-9 w=210e-9 m=1 nf=1 
m4 net5 i2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m5 net33 i1 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m6 net13 s0 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m7 net9 s1 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m8 net5 s1 net79 vss nch_hvt l=60e-9 w=320e-9 m=1 nf=1 
m9 z net79 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m10 z net79 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m11 net25 s1 net79 vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
m12 net33 i1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m13 net9 s1 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
m14 net5 i2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m15 net33 net13 net25 vdd pch_hvt l=60e-9 w=350e-9 m=1 nf=1 
m16 net13 s0 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
m17 net5 net9 net79 vdd pch_hvt l=60e-9 w=440e-9 m=1 nf=1 
m18 net37 i0 vdd vdd pch_hvt l=60e-9 w=340e-9 m=1 nf=1 
m19 net37 s0 net25 vdd pch_hvt l=60e-9 w=410e-9 m=1 nf=1 
.ends MUX3D1HVT
** End of subcircuit definition.

** Library name: civic
** Cell name: PWR_BANK
** View name: schematic
.subckt PWR_BANK code<5> code<4> code<3> code<2> code<1> code<0> dout<0> dout<1> dout<2> dout<3> dout<4> dout<5> dout<6> dout<7> dout<8> dout<9> dout<10> dout<11> dout<12> dout<13> dout<14> dout<15> en mclk rs_rising sel<1> sel<0> sysclk vdd vout vss
xi30 code<5> code<4> code<3> code<2> code<1> code<0> en ro<0> ro<64> ro<63> ro<62> ro<61> ro<60> ro<59> ro<58> ro<57> ro<56> ro<55> ro<54> ro<53> ro<52> ro<51> ro<50> ro<49> ro<48> ro<47> ro<46> ro<45> ro<44> ro<43> ro<42> ro<41> ro<40> ro<39> ro<38> ro<37> ro<36> ro<35> ro<34> ro<33> ro<32> ro<31> ro<30> ro<29> ro<28> ro<27> ro<26> ro<25> ro<24> ro<23> ro<22> ro<21> ro<20> ro<19> ro<18> ro<17> ro<16> ro<15> ro<14> ro<13> ro<12> ro<11> ro<10> ro<9> ro<8> ro<7> ro<6> ro<5> ro<4> ro<3> ro<2> ro<1> rs_rising vdd vout vss ULDO_BANK
xi16 ro<4> ro<8> ro<12> ro<16> ro<20> ro<24> ro<28> ro<32> ro<36> ro<40> ro<44> ro<48> ro<52> ro<56> ro<60> ro<64> dout<0> dout<1> dout<2> dout<3> dout<4> dout<5> dout<6> dout<7> dout<8> dout<9> dout<10> dout<11> dout<12> dout<13> dout<14> dout<15> doutn<0> doutn<1> doutn<2> doutn<3> doutn<4> doutn<5> doutn<6> doutn<7> doutn<8> doutn<9> doutn<10> doutn<11> doutn<12> doutn<13> doutn<14> doutn<15> vdd vss Dlvlxft_16B
xi28 dout<0> mclk vdd vss CKND1HVT
xi27 sysclk doutn<7> doutn<15> sel<0> sel<1> ro<0> vdd vss MUX3D1HVT
.ends PWR_BANK
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: DCAP8HVT
** View name: schematic
.subckt DCAP8HVT vdd vss
mi4 vss net9 vss vss nch_hvt l=880e-9 w=300e-9 m=1 nf=1 
m_u2 net11 net9 vss vss nch_hvt l=60e-9 w=300e-9 m=1 nf=1 
mi3 vdd net11 vdd vdd pch_hvt l=880e-9 w=430e-9 m=1 nf=1 
m_u1 net9 net11 vdd vdd pch_hvt l=60e-9 w=390e-9 m=1 nf=1 
.ends DCAP8HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: INVD1HVT
** View name: schematic
.subckt INVD1HVT i zn vdd vss
m0 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends INVD1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: AN2D4HVT
** View name: schematic
.subckt AN2D4HVT a1 a2 z vdd vss
m0 z net5 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m1 z net5 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m2 z net5 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 z net5 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m4 net5 a1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m5 net5 a1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m6 net5 a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m7 net5 a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m8 z net5 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m9 net57 a2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m10 z net5 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m11 net44 a2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m12 z net5 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m13 net5 a1 net44 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m14 net5 a1 net57 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m15 z net5 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
.ends AN2D4HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: INVD16HVT
** View name: schematic
.subckt INVD16HVT i zn vdd vss
m0 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m1 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m2 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m4 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m5 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m6 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m7 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m8 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m9 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m10 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m11 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m12 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m13 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m14 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m15 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m16 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m17 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m18 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m19 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m20 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m21 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m22 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m23 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m24 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m25 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m26 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m27 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m28 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m29 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m30 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m31 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
.ends INVD16HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: DEL015HVT
** View name: schematic
.subckt DEL015HVT i z vdd vss
m0 z net13 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi29 net25 net9 net28 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi30 net28 net9 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi37 net17 net5 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi28 net13 net9 net25 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi35 net9 net5 net44 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 net5 i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi36 net44 net5 net17 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 z net13 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi20 net57 net9 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi23 net13 net9 net25 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 net5 i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi21 net25 net9 net57 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi32 net9 net5 net44 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi31 net44 net5 net33 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi7 net33 net5 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends DEL015HVT
** End of subcircuit definition.

** Library name: civic
** Cell name: LDO_CK_GEN
** View name: schematic
.subckt LDO_CK_GEN sel_rst sysclk vdd vss
xi19 net26 net24 vdd vss INVD1HVT
xi0 sysclk net24 net25 vdd vss AN2D4HVT
xi44 net25 sel_rst vdd vss INVD16HVT
xi4 sysclk net26 vdd vss DEL015HVT
.ends LDO_CK_GEN
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: CKND0HVT
** View name: schematic
.subckt CKND0HVT i zn vdd vss
m_u2 zn i vss vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m_u1 zn i vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
.ends CKND0HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: ND3D1HVT
** View name: schematic
.subckt ND3D1HVT a1 a2 a3 zn vdd vss
m0 net9 a2 net1 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 zn a1 net9 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 net1 a3 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m3 zn a1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m4 zn a3 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m5 zn a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends ND3D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: OAI21D1HVT
** View name: schematic
.subckt OAI21D1HVT a1 a2 b zn vdd vss
m0 net9 a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u9 zn b vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m1 zn a1 net9 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u3 zn a2 net24 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m_u4 net24 b vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m_u2 zn a1 net24 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
.ends OAI21D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: ND2D1HVT
** View name: schematic
.subckt ND2D1HVT a1 a2 zn vdd vss
m0 zn a1 net1 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 net1 a2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 zn a1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends ND2D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: CKXOR2D1HVT
** View name: schematic
.subckt CKXOR2D1HVT a1 a2 z vdd vss
m0 net27 a1 net44 vdd pch_hvt l=60e-9 w=290e-9 m=1 nf=1 
m1 z net44 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m2 net5 net27 vdd vdd pch_hvt l=60e-9 w=290e-9 m=1 nf=1 
m3 net9 a1 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
m4 net5 net9 net44 vdd pch_hvt l=60e-9 w=290e-9 m=1 nf=1 
m5 net27 a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m6 net27 net9 net44 vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m7 net5 a1 net44 vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m8 net9 a1 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m9 z net44 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m10 net27 a2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m11 net5 net27 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
.ends CKXOR2D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: INVD3HVT
** View name: schematic
.subckt INVD3HVT i zn vdd vss
m0 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 zn i vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m3 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m4 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m5 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends INVD3HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: CKND6HVT
** View name: schematic
.subckt CKND6HVT i zn vdd vss
m_u1_0 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u1_3 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u1_2 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u1_4 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u1_1 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u1_5 zn i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
di3 vss i ndio_hvt area=66e-15 pj=1.18e-6 m=1
m_u2_1 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u2_3 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u2_4 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u2_0 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u2_2 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u2_5 zn i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
.ends CKND6HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: DFCNQD1HVT
** View name: schematic
.subckt DFCNQD1HVT d cp cdn q vdd vss
mi4 net53 net5 vss vss nch_hvt l=60e-9 w=350e-9 m=1 nf=1 
m0 net81 net51 net9 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 net37 net97 vss vss nch_hvt l=60e-9 w=160e-9 m=1 nf=1 
mi29 net51 net5 net44 vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi15 net37 net63 net51 vss nch_hvt l=60e-9 w=160e-9 m=1 nf=1 
m2 net63 net5 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
mi5 net97 d net53 vss nch_hvt l=60e-9 w=350e-9 m=1 nf=1 
mi49 net20 cdn vss vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi26 net44 net81 vss vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi48 net17 net37 net20 vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m3 q net81 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m4 net9 cdn vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m5 net5 cp vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
mi47 net97 net63 net17 vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m6 net5 cp vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
m7 net63 net5 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
mi43 net101 net37 vdd vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi6 net97 d net100 vdd pch_hvt l=60e-9 w=460e-9 m=1 nf=1 
m8 q net81 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi44 net101 cdn vdd vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m9 net37 net97 vdd vdd pch_hvt l=60e-9 w=220e-9 m=1 nf=1 
m10 net81 net51 vdd vdd pch_hvt l=60e-9 w=400e-9 m=1 nf=1 
mi16 net37 net5 net51 vdd pch_hvt l=60e-9 w=245e-9 m=1 nf=1 
mi24 net72 net81 vdd vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi28 net51 net63 net72 vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi45 net97 net5 net101 vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi7 net100 net63 vdd vdd pch_hvt l=60e-9 w=460e-9 m=1 nf=1 
m11 net81 cdn vdd vdd pch_hvt l=60e-9 w=400e-9 m=1 nf=1 
.ends DFCNQD1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: CKBD1HVT
** View name: schematic
.subckt CKBD1HVT i z vdd vss
m_u15 net5 i vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
mu23 z net5 vss vss nch_hvt l=60e-9 w=310e-9 m=1 nf=1 
m_u3 net5 i vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mu21 z net5 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends CKBD1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: OAI32D1HVT
** View name: schematic
.subckt OAI32D1HVT a1 a2 a3 b1 b2 zn vdd vss
m0 net17 b1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m1 net13 a1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m2 zn b2 net17 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a3 net1 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m4 net1 a2 net13 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi1 zn a1 net25 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi3 zn a3 net25 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi2 zn a2 net25 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi0 net25 b2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m_u4 net25 b1 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
.ends OAI32D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: AOI32D1HVT
** View name: schematic
.subckt AOI32D1HVT a1 a2 a3 b1 b2 zn vdd vss
mu18 zn a3 net20 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mu19 net20 b2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mu16 zn a2 net20 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mu20 net20 b1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mu17 zn a1 net20 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m0 zn a1 net21 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 zn b1 net36 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 net36 b2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m3 net25 a3 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m4 net21 a2 net25 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
.ends AOI32D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: AOI211XD0HVT
** View name: schematic
.subckt AOI211XD0HVT a1 a2 b c zn vdd vss
m_u12 zn c vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m0 zn a1 net1 vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m_u13 zn b vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m1 net1 a2 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m2 net25 b net17 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u3 net25 a1 zn vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi0 net25 a2 zn vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 net17 c vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends AOI211XD0HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: DFCSNQD4HVT
** View name: schematic
.subckt DFCSNQD4HVT d cp cdn sdn q vdd vss
m0 net81 net83 net17 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 q net81 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 net36 cdn vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m3 net24 net81 vss vss nch_hvt l=60e-9 w=210e-9 m=1 nf=1 
mi20 net5 net67 net83 vss nch_hvt l=60e-9 w=230e-9 m=1 nf=1 
m4 net61 net63 vss vss nch_hvt l=60e-9 w=210e-9 m=1 nf=1 
mi23 net63 net67 net25 vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m5 q net81 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi22 net49 net51 net83 vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi21 net63 d net29 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m6 q net81 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m7 net51 cp vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m8 net81 net83 net36 vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
mi19 net29 net51 vss vss nch_hvt l=60e-9 w=305e-9 m=1 nf=1 
mi24 net25 net5 net1 vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m9 net49 sdn net24 vss nch_hvt l=60e-9 w=210e-9 m=1 nf=1 
m10 net17 cdn vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m11 net67 net51 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m12 q net81 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m13 net5 sdn net61 vss nch_hvt l=60e-9 w=210e-9 m=1 nf=1 
mi25 net1 cdn vss vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mi33 net49 net67 net83 vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m14 q net81 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m15 net49 sdn vdd vdd pch_hvt l=60e-9 w=350e-9 m=1 nf=1 
m16 net51 cp vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m17 q net81 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m18 net5 sdn vdd vdd pch_hvt l=60e-9 w=480e-9 m=1 nf=1 
m19 net81 cdn vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi34 net63 net51 net89 vdd pch_hvt l=60e-9 w=180e-9 m=1 nf=1 
m20 net49 net81 vdd vdd pch_hvt l=60e-9 w=350e-9 m=1 nf=1 
m21 net81 net83 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi30 net5 net51 net83 vdd pch_hvt l=60e-9 w=280e-9 m=1 nf=1 
m22 net81 cdn vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m23 q net81 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m24 q net81 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi28 net96 net67 vdd vdd pch_hvt l=60e-9 w=495e-9 m=1 nf=1 
mi35 net89 net5 vdd vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m25 net5 net63 vdd vdd pch_hvt l=60e-9 w=480e-9 m=1 nf=1 
m26 net67 net51 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi26 net63 d net96 vdd pch_hvt l=60e-9 w=495e-9 m=1 nf=1 
mi36 net89 cdn vdd vdd pch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m27 net81 net83 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends DFCSNQD4HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: NR3D0HVT
** View name: schematic
.subckt NR3D0HVT a1 a2 a3 zn vdd vss
mi3 zn a1 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
mi2 zn a2 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m_u4 zn a3 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
mi1 zn a1 net13 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m_u1 net17 a3 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
mi0 net13 a2 net17 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends NR3D0HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: OR3D1HVT
** View name: schematic
.subckt OR3D1HVT a1 a2 a3 z vdd vss
m0 net13 a1 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m1 net9 a3 net1 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m2 z net9 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 net1 a2 net13 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m4 net9 a2 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m5 net9 a1 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
m6 z net9 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m7 net9 a3 vss vss nch_hvt l=60e-9 w=195e-9 m=1 nf=1 
.ends OR3D1HVT
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: NR2D1HVT
** View name: schematic
.subckt NR2D1HVT a1 a2 zn vdd vss
m0 zn a2 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m1 zn a1 vss vss nch_hvt l=60e-9 w=390e-9 m=1 nf=1 
m2 net13 a2 vdd vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a1 net13 vdd pch_hvt l=60e-9 w=520e-9 m=1 nf=1 
.ends NR2D1HVT
** End of subcircuit definition.

** Library name: model3x
** Cell name: SEL_LOGIC_V3
** View name: schematic
.subckt SEL_LOGIC_V3 nro<2> nro<1> nro<0> sel<1> sel<0> mclk srst vdd vss
xu12 n38 n90 vdd vss INVD1HVT
xu15 sel<1> n70 vdd vss INVD1HVT
xu9 cylcnt<1> n6 vdd vss INVD1HVT
xu19 nro<1> eq_99_b_0_ vdd vss INVD1HVT
xu17 nro<2> n10 vdd vss INVD1HVT
xu4 n8 eq_99_b_9_ vdd vss INVD1HVT
xu7 srst n2 vdd vss INVD1HVT
xu20 cylcnt<0> n5 vdd vss INVD1HVT
xu3 nro<0> n11 vdd vss CKND0HVT
xu6 n11 n2 eq_99_b_9_ n20 vdd vss ND3D1HVT
xu18 eq_99_b_0_ n10 n8 n7 vdd vss OAI21D1HVT
xu21 nro<0> n8 n2 n21 vdd vss OAI21D1HVT
xu5 eq_99_b_0_ n10 n8 vdd vss ND2D1HVT
xu16 nro<1> cylcnt<0> n16 vdd vss CKXOR2D1HVT
xu23 n7 cylcnt<1> n30 vdd vss CKXOR2D1HVT
xu24 cylcnt<1> cylcnt<0> n3 vdd vss CKXOR2D1HVT
xu25 eq_99_b_0_ cylcnt<0> n4 vdd vss CKXOR2D1HVT
xcknd16hvt_g1b2i1 mclk mclk_g1b1i1 vdd vss INVD3HVT
xcknd2hvt_g1b1i1 mclk_g1b1i1 mclk_g1b2i1 vdd vss CKND6HVT
xcylcnt_reg_0_ n35 mclk_g1b2i1 srst cylcnt<0> vdd vss DFCNQD1HVT
xcylcnt_reg_1_ n3 mclk_g1b2i1 srst cylcnt<1> vdd vss DFCNQD1HVT
xu28 sel<0> n38 vdd vss CKBD1HVT
xu27 n25 n37 vdd vss CKBD1HVT
xu2 n22 n36 vdd vss CKBD1HVT
xu1 n5 n35 vdd vss CKBD1HVT
xu11 n1 nro<0> n14 n12 n90 n25 vdd vss OAI32D1HVT
xu8 n16 n6 n10 cylcnt<1> n19 n12 vdd vss OAI32D1HVT
xu10 cylcnt<0> n10 nro<1> eq_99_b_9_ n5 n19 vdd vss AOI32D1HVT
xu14 n9 n11 n70 n12 n22 vdd vss AOI211XD0HVT
xsel_reg_0_ n37 mclk_g1b2i1 n21 n20 sel<0> vdd vss DFCSNQD4HVT
xsel_reg_1_ n36 mclk_g1b2i1 n20 n21 sel<1> vdd vss DFCSNQD4HVT
xu26 n4 eq_99_b_9_ n30 n9 vdd vss NR3D0HVT
xu22 n4 eq_99_b_9_ n30 n1 vdd vss OR3D1HVT
xu13 sel<0> sel<1> n14 vdd vss NR2D1HVT
.ends SEL_LOGIC_V3
** End of subcircuit definition.

** Library name: tcbn65lphvt
** Cell name: CKBD0HVT
** View name: schematic
.subckt CKBD0HVT i z vdd vss
m_u15 net5 i vss vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
mu23 z net5 vss vss nch_hvt l=60e-9 w=150e-9 m=1 nf=1 
m_u3 net5 i vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
mu21 z net5 vdd vdd pch_hvt l=60e-9 w=260e-9 m=1 nf=1 
.ends CKBD0HVT
** End of subcircuit definition.

** Library name: civic
** Cell name: DLDO_LOOP
** View name: schematic
.subckt DLDO_LOOP code<5> code<4> code<3> code<2> code<1> code<0> dout<15> dout<14> dout<13> dout<12> dout<11> dout<10> dout<9> dout<8> dout<7> dout<6> dout<5> dout<4> dout<3> dout<2> dout<1> dout<0> ldo_en nro<2> nro<1> nro<0> sel<1> sel<0> sys_clk vdd vout vss
xpwbk2 code<5> code<4> code<3> code<2> code<1> code<0> dout<15> dout<14> dout<13> dout<12> dout<11> dout<10> dout<9> dout<8> dout<7> dout<6> dout<5> dout<4> dout<3> dout<2> dout<1> dout<0> ldo_en net24 net23 sel<1> sel<0> sys_clk vdd vout vss PWR_BANK
xi0<40> vdd vss DCAP8HVT
xi0<39> vdd vss DCAP8HVT
xi0<38> vdd vss DCAP8HVT
xi0<37> vdd vss DCAP8HVT
xi0<36> vdd vss DCAP8HVT
xi0<35> vdd vss DCAP8HVT
xi0<34> vdd vss DCAP8HVT
xi0<33> vdd vss DCAP8HVT
xi0<32> vdd vss DCAP8HVT
xi0<31> vdd vss DCAP8HVT
xi0<30> vdd vss DCAP8HVT
xi0<29> vdd vss DCAP8HVT
xi0<28> vdd vss DCAP8HVT
xi0<27> vdd vss DCAP8HVT
xi0<26> vdd vss DCAP8HVT
xi0<25> vdd vss DCAP8HVT
xi0<24> vdd vss DCAP8HVT
xi0<23> vdd vss DCAP8HVT
xi0<22> vdd vss DCAP8HVT
xi0<21> vdd vss DCAP8HVT
xi0<20> vdd vss DCAP8HVT
xi0<19> vdd vss DCAP8HVT
xi0<18> vdd vss DCAP8HVT
xi0<17> vdd vss DCAP8HVT
xi0<16> vdd vss DCAP8HVT
xi0<15> vdd vss DCAP8HVT
xi0<14> vdd vss DCAP8HVT
xi0<13> vdd vss DCAP8HVT
xi0<12> vdd vss DCAP8HVT
xi0<11> vdd vss DCAP8HVT
xi0<10> vdd vss DCAP8HVT
xi0<9> vdd vss DCAP8HVT
xi0<8> vdd vss DCAP8HVT
xi0<7> vdd vss DCAP8HVT
xi0<6> vdd vss DCAP8HVT
xi0<5> vdd vss DCAP8HVT
xi0<4> vdd vss DCAP8HVT
xi0<3> vdd vss DCAP8HVT
xi0<2> vdd vss DCAP8HVT
xi0<1> vdd vss DCAP8HVT
xi0<0> vdd vss DCAP8HVT
xckgen0 net23 sys_clk vdd vss LDO_CK_GEN
xselog1 nro<2> nro<1> n1 sel<1> sel<0> net24 net23 vdd vss SEL_LOGIC_V3
xi1 nro<0> n1 vdd vss CKBD0HVT
.ends DLDO_LOOP
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: CKND3
** View name: schematic
.subckt CKND3 i zn vdd vss
m_u1_0 zn i vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u1_2 zn i vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u1_1 zn i vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u2_1 zn i vss vss nch l=60e-9 w=310e-9 m=1 nf=1 
m_u2_0 zn i vss vss nch l=60e-9 w=310e-9 m=1 nf=1 
m_u2_2 zn i vss vss nch l=60e-9 w=310e-9 m=1 nf=1 
.ends CKND3
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: CKND2D1
** View name: schematic
.subckt CKND2D1 a1 a2 zn vdd vss
m0 zn a1 net1 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 net1 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 zn a1 vdd vdd pch l=60e-9 w=390e-9 m=1 nf=1 
m3 zn a2 vdd vdd pch l=60e-9 w=390e-9 m=1 nf=1 
.ends CKND2D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: CKND1
** View name: schematic
.subckt CKND1 i zn vdd vss
m_u2 zn i vss vss nch l=60e-9 w=310e-9 m=1 nf=1 
m_u1 zn i vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends CKND1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: ND3D1
** View name: schematic
.subckt ND3D1 a1 a2 a3 zn vdd vss
m0 net9 a2 net1 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 zn a1 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 net1 a3 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m3 zn a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m4 zn a3 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m5 zn a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends ND3D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: NR2XD0
** View name: schematic
.subckt NR2XD0 a1 a2 zn vdd vss
m0 zn a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m1 zn a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m2 net13 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a1 net13 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends NR2XD0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: MUX2ND0
** View name: schematic
.subckt MUX2ND0 i0 i1 s zn vdd vss
m0 net37 s vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi111 net13 i0 vdd vdd pch l=60e-9 w=310e-9 m=1 nf=1 
mi24 net9 i1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi5 zn s net13 vdd pch l=60e-9 w=390e-9 m=1 nf=1 
mi25 zn net37 net9 vdd pch l=60e-9 w=390e-9 m=1 nf=1 
m1 net37 s vss vss nch l=60e-9 w=210e-9 m=1 nf=1 
mi20 net33 i1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi12 zn net37 net32 vss nch l=60e-9 w=230e-9 m=1 nf=1 
mi21 zn s net33 vss nch l=60e-9 w=230e-9 m=1 nf=1 
mi19 net32 i0 vss vss nch l=60e-9 w=230e-9 m=1 nf=1 
.ends MUX2ND0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OA31D1
** View name: schematic
.subckt OA31D1 a1 a2 a3 b z vdd vss
m0 z net25 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi6 net5 a1 net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u5 vss b net5 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi8 net5 a3 net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi7 net5 a2 net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi3 net37 a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi4 net33 a2 net37 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 z net25 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u11 net25 b vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi5 net25 a3 net33 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends OA31D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: CKBD1
** View name: schematic
.subckt CKBD1 i z vdd vss
m_u15 net5 i vss vss nch l=60e-9 w=310e-9 m=1 nf=1 
mu23 z net5 vss vss nch l=60e-9 w=310e-9 m=1 nf=1 
m_u3 net5 i vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mu21 z net5 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends CKBD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: NR4D0
** View name: schematic
.subckt NR4D0 a1 a2 a3 a4 zn vdd vss
mi34 zn a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi5 zn a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi35 zn a3 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi36 zn a4 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi27 net29 a2 net32 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi28 zn a1 net29 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi26 net32 a3 net24 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi7 net24 a4 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends NR4D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: AN3XD1
** View name: schematic
.subckt AN3XD1 a1 a2 a3 z vdd vss
m0 net13 a3 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 z net11 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 net5 a2 net13 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m3 net11 a1 net5 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m4 z net11 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m5 net11 a3 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m6 net11 a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m7 net11 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends AN3XD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OA211D1
** View name: schematic
.subckt OA211D1 a1 a2 b c z vdd vss
mi17 net17 c vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi15 net25 a1 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi16 net9 b net17 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m0 z net25 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi7 net25 a2 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi13 net37 a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi12 net25 c vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u12 net25 b vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi14 net25 a2 net37 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 z net25 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends OA211D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: DFCSNQD1
** View name: schematic
.subckt DFCSNQD1 d cp cdn sdn q vdd vss
m0 net61 net100 net37 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 q net61 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 net20 net61 vss vss nch l=60e-9 w=210e-9 m=1 nf=1 
mi20 net97 net81 net100 vss nch l=60e-9 w=230e-9 m=1 nf=1 
m3 net45 net47 vss vss nch l=60e-9 w=210e-9 m=1 nf=1 
mi23 net47 net81 net44 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m4 net37 cdn vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi22 net125 net13 net100 vss nch l=60e-9 w=150e-9 m=1 nf=1 
mi21 net47 d net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi19 net25 net13 vss vss nch l=60e-9 w=305e-9 m=1 nf=1 
mi24 net44 net97 net5 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m5 net125 sdn net20 vss nch l=60e-9 w=210e-9 m=1 nf=1 
m6 net13 cp vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m7 net97 sdn net45 vss nch l=60e-9 w=210e-9 m=1 nf=1 
mi25 net5 cdn vss vss nch l=60e-9 w=150e-9 m=1 nf=1 
m8 net81 net13 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi33 net125 net81 net100 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
m9 net125 sdn vdd vdd pch l=60e-9 w=350e-9 m=1 nf=1 
m10 net61 net100 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m11 q net61 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m12 net97 sdn vdd vdd pch l=60e-9 w=480e-9 m=1 nf=1 
mi34 net47 net13 net108 vdd pch l=60e-9 w=180e-9 m=1 nf=1 
m13 net125 net61 vdd vdd pch l=60e-9 w=350e-9 m=1 nf=1 
mi30 net97 net13 net100 vdd pch l=60e-9 w=280e-9 m=1 nf=1 
m14 net61 cdn vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m15 net13 cp vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi28 net72 net81 vdd vdd pch l=60e-9 w=495e-9 m=1 nf=1 
m16 net81 net13 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi35 net108 net97 vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
m17 net97 net47 vdd vdd pch l=60e-9 w=480e-9 m=1 nf=1 
mi26 net47 d net72 vdd pch l=60e-9 w=495e-9 m=1 nf=1 
mi36 net108 cdn vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
.ends DFCSNQD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: AOI21D1
** View name: schematic
.subckt AOI21D1 a1 a2 b zn vdd vss
m_u3 net5 a1 zn vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u2 net5 b vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u4 net5 a2 zn vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi2 zn a1 net13 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u7 zn b vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi3 net13 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
.ends AOI21D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: AO221D0
** View name: schematic
.subckt AO221D0 a1 a2 b1 b2 c z vdd vss
mu22 vdd c net9 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi9 net13 a2 net20 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi10 net13 a1 net20 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi6 net9 b2 net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m0 z net20 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi7 net9 b1 net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m1 net20 a1 net33 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m2 net20 b1 net25 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m3 z net20 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m4 net33 a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mu20 net20 c vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m5 net25 b2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends AO221D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OAI211D1
** View name: schematic
.subckt OAI211D1 a1 a2 b c zn vdd vss
mi3 net13 c vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi2 net9 b net13 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u3 zn a2 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u2 zn a1 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi1 zn a2 net25 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi0 net25 a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u11 zn c vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u12 zn b vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends OAI211D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: ND2D1
** View name: schematic
.subckt ND2D1 a1 a2 zn vdd vss
m0 zn a1 net1 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 net1 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 zn a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends ND2D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: MUX3ND0
** View name: schematic
.subckt MUX3ND0 i0 i1 i2 s0 s1 zn vdd vss
m0 net25 s0 net20 vdd pch l=60e-9 w=410e-9 m=1 nf=1 
m1 net29 i2 vdd vdd pch l=60e-9 w=540e-9 m=1 nf=1 
m2 net25 i0 vdd vdd pch l=60e-9 w=310e-9 m=1 nf=1 
m3 net51 s1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m4 net5 net13 net20 vdd pch l=60e-9 w=360e-9 m=1 nf=1 
m5 net13 s0 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m6 net20 s1 zn vdd pch l=60e-9 w=280e-9 m=1 nf=1 
m7 net5 i1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m8 net29 net51 zn vdd pch l=60e-9 w=280e-9 m=1 nf=1 
m9 net5 s0 net20 vss nch l=60e-9 w=240e-9 m=1 nf=1 
m10 net25 i0 vss vss nch l=60e-9 w=230e-9 m=1 nf=1 
m11 net5 i1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m12 net29 s1 zn vss nch l=60e-9 w=210e-9 m=1 nf=1 
m13 net13 s0 vss vss nch l=60e-9 w=210e-9 m=1 nf=1 
m14 net20 net51 zn vss nch l=60e-9 w=210e-9 m=1 nf=1 
m15 net25 net13 net20 vss nch l=60e-9 w=260e-9 m=1 nf=1 
m16 net29 i2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m17 net51 s1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
.ends MUX3ND0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OAI22D1
** View name: schematic
.subckt OAI22D1 a1 a2 b1 b2 zn vdd vss
m_u3 zn a1 net5 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u5 net5 b1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u4 net5 b2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u2 zn a2 net5 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi1 zn b1 net32 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi3 zn a1 net17 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mu24 net32 b2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi2 net17 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends OAI22D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: HA1D0
** View name: schematic
.subckt HA1D0 a b s co vdd vss
m0 net9 a vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 net13 net5 net72 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m2 net25 a vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m3 co net25 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m4 net25 b vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m5 net13 net9 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m6 net9 b net72 vdd pch l=60e-9 w=310e-9 m=1 nf=1 
m7 net5 b vdd vdd pch l=60e-9 w=285e-9 m=1 nf=1 
m8 s net72 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m9 net9 net5 net72 vss nch l=60e-9 w=205e-9 m=1 nf=1 
m10 net56 b vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m11 net9 a vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m12 s net72 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m13 net25 a net56 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m14 net13 b net72 vss nch l=60e-9 w=290e-9 m=1 nf=1 
m15 net5 b vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m16 net13 net9 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m17 co net25 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends HA1D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: CKXOR2D1
** View name: schematic
.subckt CKXOR2D1 a1 a2 z vdd vss
m0 net27 a1 net44 vdd pch l=60e-9 w=290e-9 m=1 nf=1 
m1 z net44 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m2 net5 net27 vdd vdd pch l=60e-9 w=290e-9 m=1 nf=1 
m3 net9 a1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m4 net5 net9 net44 vdd pch l=60e-9 w=290e-9 m=1 nf=1 
m5 net27 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m6 net27 net9 net44 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m7 net5 a1 net44 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m8 net9 a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m9 z net44 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m10 net27 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m11 net5 net27 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends CKXOR2D1
** End of subcircuit definition.

** Library name: civicR
** Cell name: DLDO_LOGIC_V1_DW01_inc_0
** View name: schematic
.subckt DLDO_LOGIC_V1_DW01_inc_0 sum<6> sum<5> sum<4> sum<3> sum<2> sum<1> sum<0> a<6> a<5> a<4> a<3> a<2> a<1> a<0> vss vdd
xu2 a<0> sum<0> vdd vss INVD1
xu1_1_5 a<5> carry<5> sum<5> carry<6> vdd vss HA1D0
xu1_1_3 a<3> carry<3> sum<3> carry<4> vdd vss HA1D0
xu1_1_4 a<4> carry<4> sum<4> carry<5> vdd vss HA1D0
xu1_1_2 a<2> carry<2> sum<2> carry<3> vdd vss HA1D0
xu1_1_1 a<1> a<0> sum<1> carry<2> vdd vss HA1D0
xu1 carry<6> a<6> sum<6> vdd vss CKXOR2D1
.ends DLDO_LOGIC_V1_DW01_inc_0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: AO21D1
** View name: schematic
.subckt AO21D1 a1 a2 b z vdd vss
m_u7 net5 a1 net1 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m0 z net5 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi6 net5 b vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi7 net1 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u3 net25 a1 net5 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u2 net25 b vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m_u4 net25 a2 net5 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 z net5 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends AO21D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: XNR2D1
** View name: schematic
.subckt XNR2D1 a1 a2 zn vdd vss
m0 net27 net9 net44 vdd pch l=60e-9 w=370e-9 m=1 nf=1 
m1 zn net44 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m2 net5 net27 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m3 net9 a1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m4 net5 a1 net44 vdd pch l=60e-9 w=235e-9 m=1 nf=1 
m5 net27 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m6 net27 a1 net44 vss nch l=60e-9 w=225e-9 m=1 nf=1 
m7 net5 net9 net44 vss nch l=60e-9 w=190e-9 m=1 nf=1 
m8 net9 a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m9 zn net44 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m10 net27 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m11 net5 net27 vss vss nch l=60e-9 w=190e-9 m=1 nf=1 
.ends XNR2D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: ND4D1
** View name: schematic
.subckt ND4D1 a1 a2 a3 a4 zn vdd vss
mi3 net13 a2 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi4 net9 a3 net1 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mu53 zn a1 net13 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi5 net1 a4 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi1 zn a3 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi2 zn a4 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi0 zn a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi7 zn a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends ND4D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: INR3D0
** View name: schematic
.subckt INR3D0 a1 b1 b2 zn vdd vss
m0 net13 net9 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 net9 a1 vdd vdd pch l=60e-9 w=270e-9 m=1 nf=1 
m2 zn b2 net1 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m3 net1 b1 net13 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m4 zn b2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m5 zn net9 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m6 zn b1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m7 net9 a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends INR3D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: AN2XD1
** View name: schematic
.subckt AN2XD1 a1 a2 z vdd vss
m0 net9 a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 net5 a1 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 z net5 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m3 z net5 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m4 net5 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m5 net5 a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends AN2XD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: NR2D1
** View name: schematic
.subckt NR2D1 a1 a2 zn vdd vss
m0 zn a2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 zn a1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 net13 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a1 net13 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends NR2D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: MAOI222D1
** View name: schematic
.subckt MAOI222D1 a b c zn vdd vss
mi1 net5 b zn vss nch l=60e-9 w=210e-9 m=1 nf=1 
mi4 net13 b vss vss nch l=60e-9 w=210e-9 m=1 nf=1 
mu6 zn a net13 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mu9 net5 a zn vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi5 net5 c vss vss nch l=60e-9 w=210e-9 m=1 nf=1 
mu5 net33 a zn vdd pch l=60e-9 w=455e-9 m=1 nf=1 
mu4 net33 b zn vdd pch l=60e-9 w=455e-9 m=1 nf=1 
mi3 net33 c vdd vdd pch l=60e-9 w=455e-9 m=1 nf=1 
mi2 zn a net28 vdd pch l=60e-9 w=455e-9 m=1 nf=1 
mu2 net28 b vdd vdd pch l=60e-9 w=455e-9 m=1 nf=1 
.ends MAOI222D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: MOAI22D1
** View name: schematic
.subckt MOAI22D1 a1 a2 b1 b2 zn vdd vss
mu1 net37 b1 net20 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi6 net9 net37 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mu9 net9 a1 zn vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi5 net20 b2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mu10 net9 a2 zn vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi1 net37 b1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi3 net33 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi4 zn a1 net33 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi2 zn net37 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mu3 net37 b2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends MOAI22D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OA32D0
** View name: schematic
.subckt OA32D0 a1 a2 a3 b1 b2 z vdd vss
m0 z net5 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m1 net17 b1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m2 net13 a1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m3 net5 b2 net17 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m4 net5 a3 net1 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m5 net1 a2 net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi3 net5 a3 net33 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m6 z net5 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi11 net33 b2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi12 net33 b1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi8 net5 a2 net33 vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi9 net5 a1 net33 vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends OA32D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: IOA21D1
** View name: schematic
.subckt IOA21D1 a1 a2 b zn vdd vss
m0 net5 a2 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m1 zn b vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m2 net5 a1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m3 zn net5 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m4 net29 a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m5 net5 a1 net29 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m6 zn b net24 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m7 net24 net5 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
.ends IOA21D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OAI32D1
** View name: schematic
.subckt OAI32D1 a1 a2 a3 b1 b2 zn vdd vss
m0 net17 b1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 net13 a1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m2 zn b2 net17 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m3 zn a3 net1 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m4 net1 a2 net13 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi1 zn a1 net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi3 zn a3 net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi2 zn a2 net25 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi0 net25 b2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m_u4 net25 b1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
.ends OAI32D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OR2D1
** View name: schematic
.subckt OR2D1 a1 a2 z vdd vss
m0 z net5 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 net5 a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m2 net5 a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m3 z net5 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m4 net17 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m5 net5 a1 net17 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends OR2D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: INR2D1
** View name: schematic
.subckt INR2D1 a1 b1 zn vdd vss
m0 zn net11 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 zn b1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 net11 a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m3 net11 a1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m4 zn b1 net20 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m5 net20 net11 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends INR2D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: AOI221D0
** View name: schematic
.subckt AOI221D0 a1 a2 b1 b2 c zn vdd vss
mu22 vdd c net20 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi9 net13 a1 zn vdd pch l=60e-9 w=280e-9 m=1 nf=1 
mi6 net20 b2 net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi7 net20 b1 net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi8 net13 a2 zn vdd pch l=60e-9 w=280e-9 m=1 nf=1 
m0 zn b1 net29 vss nch l=60e-9 w=195e-9 m=1 nf=1 
mu20 zn c vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m1 net29 b2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m2 zn a1 net28 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m3 net28 a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends AOI221D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OA22D0
** View name: schematic
.subckt OA22D0 a1 a2 b1 b2 z vdd vss
m0 z net5 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi18 net13 b1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi20 net5 a1 net13 vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi19 net5 a2 net13 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m_u4 net13 b2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m1 z net5 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mu24 net33 b2 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi17 net5 a1 net32 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi15 net5 b1 net33 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi16 net32 a2 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
.ends OA22D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: MUX2D0
** View name: schematic
.subckt MUX2D0 i0 i1 s z vdd vss
m0 z net5 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m1 net17 s vdd vdd pch l=60e-9 w=250e-9 m=1 nf=1 
mi111 net13 i0 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi24 net9 i1 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi5 net5 s net13 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi25 net5 net17 net9 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m2 net17 s vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi20 net36 i1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi12 net5 net17 net25 vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi21 net5 s net36 vss nch l=60e-9 w=195e-9 m=1 nf=1 
m3 z net5 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi19 net25 i0 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
.ends MUX2D0
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: DFCNQD1
** View name: schematic
.subckt DFCNQD1 d cp cdn q vdd vss
mi4 net53 net5 vss vss nch l=60e-9 w=350e-9 m=1 nf=1 
m0 net81 net51 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 net37 net97 vss vss nch l=60e-9 w=160e-9 m=1 nf=1 
mi29 net51 net5 net44 vss nch l=60e-9 w=150e-9 m=1 nf=1 
mi15 net37 net63 net51 vss nch l=60e-9 w=160e-9 m=1 nf=1 
m2 net63 net5 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi5 net97 d net53 vss nch l=60e-9 w=350e-9 m=1 nf=1 
mi49 net20 cdn vss vss nch l=60e-9 w=150e-9 m=1 nf=1 
mi26 net44 net81 vss vss nch l=60e-9 w=150e-9 m=1 nf=1 
mi48 net17 net37 net20 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m3 q net81 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m4 net9 cdn vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m5 net5 cp vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi47 net97 net63 net17 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m6 net5 cp vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m7 net63 net5 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi43 net101 net37 vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi6 net97 d net100 vdd pch l=60e-9 w=460e-9 m=1 nf=1 
m8 q net81 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi44 net101 cdn vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
m9 net37 net97 vdd vdd pch l=60e-9 w=220e-9 m=1 nf=1 
m10 net81 net51 vdd vdd pch l=60e-9 w=400e-9 m=1 nf=1 
mi16 net37 net5 net51 vdd pch l=60e-9 w=245e-9 m=1 nf=1 
mi24 net72 net81 vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi28 net51 net63 net72 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi45 net97 net5 net101 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi7 net100 net63 vdd vdd pch l=60e-9 w=460e-9 m=1 nf=1 
m11 net81 cdn vdd vdd pch l=60e-9 w=400e-9 m=1 nf=1 
.ends DFCNQD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: DFD1
** View name: schematic
.subckt DFD1 d cp q qn vdd vss
m0 net67 net100 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m1 qn net97 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi4 net20 net13 vss vss nch l=60e-9 w=370e-9 m=1 nf=1 
mi55 net97 net13 net100 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m2 net11 net17 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi50 net11 net99 net100 vss nch l=60e-9 w=200e-9 m=1 nf=1 
m3 net97 net67 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m4 net99 net13 vss vss nch l=60e-9 w=180e-9 m=1 nf=1 
mi5 net17 d net20 vss nch l=60e-9 w=370e-9 m=1 nf=1 
m5 net13 cp vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
mi48 net9 net11 vss vss nch l=60e-9 w=150e-9 m=1 nf=1 
m6 q net67 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi47 net17 net99 net9 vss nch l=60e-9 w=150e-9 m=1 nf=1 
m7 net67 net100 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi54 net97 net99 net100 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
m8 net99 net13 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi43 net60 net11 vdd vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi6 net17 d net53 vdd pch l=60e-9 w=460e-9 m=1 nf=1 
m9 qn net97 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m10 net13 cp vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m11 q net67 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m12 net11 net17 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m13 net97 net67 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
mi52 net11 net13 net100 vdd pch l=60e-9 w=215e-9 m=1 nf=1 
mi45 net17 net13 net60 vdd pch l=60e-9 w=150e-9 m=1 nf=1 
mi7 net53 net99 vdd vdd pch l=60e-9 w=460e-9 m=1 nf=1 
.ends DFD1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: OA222D1
** View name: schematic
.subckt OA222D1 a1 a2 b1 b2 c1 c2 z vdd vss
mu25 net9 c1 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi18 net33 a2 net20 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi17 net33 a1 net20 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi15 net20 b1 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi14 net9 c2 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi16 net20 b2 net9 vss nch l=60e-9 w=390e-9 m=1 nf=1 
m0 z net33 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
mi13 net33 a1 net56 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi2 net49 c1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi11 net45 b1 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi12 net56 a2 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m1 z net33 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi8 net33 c2 net49 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
mi9 net33 b2 net45 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
.ends OA222D1
** End of subcircuit definition.

** Library name: tcbn65lp
** Cell name: IAO21D1
** View name: schematic
.subckt IAO21D1 a1 a2 b zn vdd vss
m0 net11 a2 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m1 zn net11 vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m2 zn b vss vss nch l=60e-9 w=390e-9 m=1 nf=1 
m3 net11 a1 vss vss nch l=60e-9 w=195e-9 m=1 nf=1 
m4 zn b net25 vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m5 net25 net11 vdd vdd pch l=60e-9 w=520e-9 m=1 nf=1 
m6 net11 a1 net24 vdd pch l=60e-9 w=260e-9 m=1 nf=1 
m7 net24 a2 vdd vdd pch l=60e-9 w=260e-9 m=1 nf=1 
.ends IAO21D1
** End of subcircuit definition.

** Library name: civicR
** Cell name: DLDO_LOGIC_V1
** View name: schematic
.subckt DLDO_LOGIC_V1 thm2bin<4> thm2bin<3> thm2bin<2> thm2bin<1> thm2bin<0> clk en_ldo boost mode code<5> code<4> code<3> code<2> code<1> code<0> cfg_2<5> cfg_2<4> cfg_2<3> cfg_2<2> cfg_2<1> cfg_2<0> din<15> din<14> din<13> din<12> din<11> din<10> din<9> din<8> din<7> din<6> din<5> din<4> din<3> din<2> din<1> din<0> cfg_1<5> cfg_1<4> cfg_1<3> cfg_1<2> cfg_1<1> cfg_1<0> sel<1> sel<0> vdd vss
xu123 n935 n157 n45 vdd vss CKND2D1
xu124 cfg_2<5> n157 n140 vdd vss CKND2D1
xu155 n941 n940 n942 vdd vss CKND2D1
xu115 cfg_2<4> n157 n139 vdd vss CKND2D1
xu114 n927 n157 n44 vdd vss CKND2D1
xu47 n52 n1 n930 vdd vss CKND2D1
xu51 n936 n894 n896 vdd vss CKND2D1
xu103 cfg_2<0> n157 n179 vdd vss CKND2D1
xu102 n917 n157 n178 vdd vss CKND2D1
xu76 n903 n1 n907 vdd vss CKND2D1
xu110 n157 cfg_2<1> n181 vdd vss CKND2D1
xu109 n157 n922 n180 vdd vss CKND2D1
xu99 cfg_2<3> n157 n138 vdd vss CKND2D1
xu97 n915 n157 n43 vdd vss CKND2D1
xu80 n157 cfg_2<2> n137 vdd vss CKND2D1
xu79 n157 n906 n46 vdd vss CKND2D1
xu87 n908 n907 n909 vdd vss CKND2D1
xu170 n951 n950 n381 vdd vss CKND2D1
xu67 n177 n900 n918 vdd vss CKND2D1
xu168 n951 n949 code<4> vdd vss CKND2D1
xu166 n951 n948 code<3> vdd vss CKND2D1
xu164 n951 n947 code<2> vdd vss CKND2D1
xu162 n951 n946 code<1> vdd vss CKND2D1
xu160 n951 n945 code<0> vdd vss CKND2D1
xu57 n889 n952 n57 vdd vss CKND2D1
xu158 mode code_reg<6> n951 vdd vss CKND2D1
xu118 n937 n928 vdd vss CKND1
xu116 code_reg<4> n929 vdd vss CKND1
xu172 cfg_1<0> n957 vdd vss CKND1
xu122 cfg_2<5> n935 vdd vss CKND1
xu60 n27 n938 vdd vss CKND1
xu113 cfg_2<4> n927 vdd vss CKND1
xu50 code_reg<6> n894 vdd vss CKND1
xu171 cfg_1<1> n956 vdd vss CKND1
xu173 cfg_1<2> n955 vdd vss CKND1
xu174 cfg_1<3> n954 vdd vss CKND1
xu49 code_reg<5> n936 vdd vss CKND1
xu2 n930 n2 vdd vss CKND1
xu74 n54 n901 vdd vss CKND1
xu78 cfg_2<2> n906 vdd vss CKND1
xu58 n57 n899 vdd vss CKND1
xu59 n177 n898 vdd vss CKND1
xu45 n62 n952 vdd vss CKND1
xu66 n58 n900 vdd vss CKND1
xu56 n52 n895 vdd vss CKND1
xu100 cfg_2<0> n917 vdd vss CKND1
xu1 boost n1 vdd vss CKND1
xu68 n918 n924 vdd vss CKND1
xu104 cfg_2<1> n922 vdd vss CKND1
xu84 cfg_2<3> n915 vdd vss CKND1
xu54 code_reg<1> n897 vdd vss CKND1
xu53 code_reg<3> n911 vdd vss CKND1
xu52 code_reg<2> n912 vdd vss CKND1
xu117 code_reg<4> n890 n2 n937 vdd vss ND3D1
xu65 n63 n62 n889 n58 vdd vss ND3D1
xu55 n912 n911 n897 n923 vdd vss ND3D1
xu153 n937 n936 n943 vdd vss NR2XD0
xu69 n52 n924 n902 vdd vss NR2XD0
xu105 boost n918 n919 vdd vss NR2XD0
xu111 n924 n923 n925 vdd vss NR2XD0
xu121 n933 n941 code_reg<5> n934 vdd vss MUX2ND0
xu154 n2 n938 code_reg<5> n940 vdd vss MUX2ND0
xu156 n943 n942 code_reg<6> n944 vdd vss MUX2ND0
xu120 n930 n27 code_reg<4> n932 vdd vss MUX2ND0
xu75 n902 n901 code_reg<1> n903 vdd vss MUX2ND0
xu106 n2 n919 code_reg<1> n921 vdd vss MUX2ND0
xu77 n904 n907 code_reg<2> n905 vdd vss MUX2ND0
xu86 n2 n938 code_reg<2> n908 vdd vss MUX2ND0
xu90 n910 n909 code_reg<3> n914 vdd vss MUX2ND0
xu169 cfg_1<5> code_reg<5> mode n950 vdd vss MUX2ND0
xu167 cfg_1<4> code_reg<4> mode n949 vdd vss MUX2ND0
xu165 cfg_1<3> code_reg<3> mode n948 vdd vss MUX2ND0
xu163 cfg_1<2> code_reg<2> mode n947 vdd vss MUX2ND0
xu161 cfg_1<1> code_reg<1> mode n946 vdd vss MUX2ND0
xu159 cfg_1<0> n177 mode n945 vdd vss MUX2ND0
xu7 n896 code_reg<4> n923 n895 n889 vdd vss OA31D1
xu44 n381 code<5> vdd vss CKBD1
xu4 boost n952 n63 n52 n886 vdd vss NR4D0
xu8 code_reg<3> code_reg<1> code_reg<2> n890 vdd vss AN3XD1
xu5 n888 n912 n911 n887 vdd vss AN3XD1
xu85 code_reg<2> code_reg<1> n2 n910 vdd vss AN3XD1
xu6 n899 n898 n938 n897 n888 vdd vss OA211D1
xcode_reg_reg_5_ n136 clk n45 n140 code_reg<5> vdd vss DFCSNQD1
xcode_reg_reg_4_ n230 clk n44 n139 code_reg<4> vdd vss DFCSNQD1
xcode_reg_reg_0_ n226 clk n178 n179 n177 vdd vss DFCSNQD1
xcode_reg_reg_1_ n227 clk n180 n181 code_reg<1> vdd vss DFCSNQD1
xcode_reg_reg_3_ n229 clk n43 n138 code_reg<3> vdd vss DFCSNQD1
xcode_reg_reg_2_ n228 clk n46 n137 code_reg<2> vdd vss DFCSNQD1
xu119 n887 n929 n928 n933 vdd vss AOI21D1
xu15 n79 n109 n80 n106 vdd vss AOI21D1
xu21 din<15> din<9> n112 n111 vdd vss AOI21D1
xu107 n203 n886 n888 n920 vdd vss AOI21D1
xu91 n205 n886 n887 n913 vdd vss AOI21D1
xu64 n2 code_reg<1> n888 n904 vdd vss AOI21D1
xu3 n206 n886 cfg_2<4> boost n926 n230 vdd vss AO221D0
xu31 n207 n886 cfg_2<5> boost n934 n136 vdd vss AO221D0
xu32 n177 n2 n202 n886 n916 n226 vdd vss AO221D0
xu28 n204 n886 cfg_2<2> boost n905 n228 vdd vss AO221D0
xu108 n1 n922 n921 n920 n227 vdd vss OAI211D1
xu95 n1 n915 n914 n913 n229 vdd vss OAI211D1
xu11 n65 n734 n71 vdd vss ND2D1
xu14 n54 n1 n27 vdd vss ND2D1
xu10 n58 n57 n54 vdd vss ND2D1
xu101 n58 n57 n917 n177 boost n916 vdd vss MUX3ND0
xu22 din<1> n15 din<3> n78 n791 vdd vss OAI22D1
xu20 din<13> n76 din<7> n77 n777 vdd vss OAI22D1
xu27 din<0> n81 din<10> n82 n768 vdd vss OAI22D1
xu112 n27 n925 n890 n930 n931 vdd vss OAI22D1
xadd_46 n208 n207 n206 n205 n204 n203 n202 code_reg<6> code_reg<5> code_reg<4> code_reg<3> code_reg<2> code_reg<1> n177 vss vdd DLDO_LOGIC_V1_DW01_inc_0
xu139 n105 n103 n116 vdd vss CKXOR2D1
xu138 n94 n93 n779 vdd vss CKXOR2D1
xu136 n777 n112 n94 vdd vss CKXOR2D1
xu137 n110 n95 n93 vdd vss CKXOR2D1
xu135 n733 n791 n95 vdd vss CKXOR2D1
xu150 n88 n87 n108 vdd vss CKXOR2D1
xu148 din<13> din<12> n88 vdd vss CKXOR2D1
xu149 din<7> din<2> n87 vdd vss CKXOR2D1
xu134 n97 n96 n741 vdd vss CKXOR2D1
xu132 n768 n113 n97 vdd vss CKXOR2D1
xu133 n109 n98 n96 vdd vss CKXOR2D1
xu131 n731 n767 n98 vdd vss CKXOR2D1
xu146 n90 n89 n114 vdd vss CKXOR2D1
xu144 din<10> din<8> n90 vdd vss CKXOR2D1
xu145 din<4> din<0> n89 vdd vss CKXOR2D1
xu143 n92 n91 n107 vdd vss CKXOR2D1
xu141 din<14> din<11> n92 vdd vss CKXOR2D1
xu142 din<6> din<5> n91 vdd vss CKXOR2D1
xu63 n70 n71 n885 vdd vss CKXOR2D1
xu128 n101 n100 n18 vdd vss CKXOR2D1
xu126 n728 n732 n101 vdd vss CKXOR2D1
xu127 n106 n102 n100 vdd vss CKXOR2D1
xu125 n739 n734 n102 vdd vss CKXOR2D1
xu130 n741 n99 n115 vdd vss CKXOR2D1
xu129 n104 n779 n99 vdd vss CKXOR2D1
xu152 n111 n86 n736 vdd vss CKXOR2D1
xu151 din<3> din<1> n86 vdd vss CKXOR2D1
xu147 n736 n108 n105 vdd vss CKXOR2D1
xu140 n114 n107 n103 vdd vss CKXOR2D1
xu93 n731 n767 n79 vdd vss CKXOR2D1
xu73 n791 n112 n74 vdd vss CKXOR2D1
xu96 din<6> din<14> n84 vdd vss CKXOR2D1
xu23 n111 n15 vdd vss INVD1
xu9 n739 n14 vdd vss INVD1
xu37 din<11> n17 vdd vss INVD1
xu30 n2 n890 n887 n891 vdd vss AO21D1
xu62 n956 n115 n116 n69 vdd vss AO21D1
xu89 din<4> din<8> n113 n81 vdd vss AO21D1
xu71 din<2> din<12> n76 vdd vss XNR2D1
xu83 n106 n734 n72 vdd vss XNR2D1
xu19 n65 n732 n66 n734 n62 vdd vss ND4D1
xu41 n113 din<0> din<10> n65 vdd vss INR3D0
xu40 n731 din<11> din<5> n734 vdd vss INR3D0
xu38 n112 din<1> din<3> n732 vdd vss INR3D0
xu39 n733 din<13> din<7> n66 vdd vss INR3D0
xu70 n76 din<13> n77 vdd vss AN2XD1
xu88 n81 din<0> n82 vdd vss AN2XD1
xu82 n105 n103 n104 vdd vss AN2XD1
xu72 n108 n736 n110 vdd vss AN2XD1
xu92 n114 n107 n109 vdd vss AN2XD1
xu36 n84 n17 n83 vdd vss NR2D1
xu33 n932 n931 n941 vdd vss NR2D1
xu25 din<9> din<15> n112 vdd vss NR2D1
xu42 din<12> din<2> n733 vdd vss NR2D1
xu26 din<4> din<8> n113 vdd vss NR2D1
xu43 din<14> din<6> n731 vdd vss NR2D1
xu81 n779 n104 n741 n739 vdd vss MAOI222D1
xu94 din<5> n83 n17 n84 n767 vdd vss MOAI22D1
xu16 n79 n109 n65 n113 n768 n80 vdd vss OA32D0
xu157 n208 n886 n944 n377 vdd vss IOA21D1
xu17 n74 n110 n75 n728 vdd vss IOA21D1
xu18 n74 n110 n66 n777 n733 n75 vdd vss OAI32D1
xu98 sel<0> sel<1> n52 vdd vss OR2D1
xu24 din<1> n111 n78 vdd vss INR2D1
xu35 n954 n885 n955 n18 n68 n892 vdd vss AOI221D0
xu12 n72 n14 n732 n66 n73 n70 vdd vss AOI221D0
xu13 n72 n14 n728 n732 n73 vdd vss OA22D0
xu29 n891 n931 code_reg<4> n926 vdd vss MUX2D0
xcode_reg_reg_6_ n377 clk en_ldo_reg code_reg<6> vdd vss DFCNQD1
xen_ldo_reg_reg en_ldo clk en_ldo_reg n157 vdd vss DFD1
xu61 n115 n956 n957 n69 n18 n955 n68 vdd vss OA222D1
xu34 n885 n954 n892 n63 vdd vss IAO21D1
.ends DLDO_LOGIC_V1
** End of subcircuit definition.

** Library name: civicR
** Cell name: DLDO_TOP
** View name: schematic
xi5 ldo_en sys_clk net012 vdd vss DFQD1
xi3 net012 net014 vdd vss INVD1
xloop0 code<5> code<4> code<3> code<2> code<1> code<0> net22<0> net22<1> net22<2> net22<3> net22<4> net22<5> net22<6> net22<7> net22<8> net22<9> net22<10> net22<11> net22<12> net22<13> net22<14> net22<15> net011 nro<2> nro<1> nro<0> sel<1> sel<0> sys_clk_cts_0 vdd vout vss DLDO_LOOP
xi4 net014 net011 vdd vss CKND3
xlogic1 net23<0> net23<1> net23<2> net23<3> net23<4> sys_clk net011 boost mode code<5> code<4> code<3> code<2> code<1> code<0> cfg_2<5> cfg_2<4> cfg_2<3> cfg_2<2> cfg_2<1> cfg_2<0> net22<0> net22<1> net22<2> net22<3> net22<4> net22<5> net22<6> net22<7> net22<8> net22<9> net22<10> net22<11> net22<12> net22<13> net22<14> net22<15> cfg_1<5> cfg_1<4> cfg_1<3> cfg_1<2> cfg_1<1> cfg_1<0> sel<1> sel<0> vdd vss DLDO_LOGIC_V1
.END
